`timescale 1ns / 1ps

module CBTest(
    
    );
endmodule
