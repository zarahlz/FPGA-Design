module t();
    wire a;
    wire b;

    assign a = b;
    assign b = a;

endmodule